`timescale 1ns / 1ps

module storage(
    );


endmodule
